package PCIe_pkg;
  
    import uvm_pkg::*;
    
    `include "Defines.sv"
    `include "uvm_macros.svh"
    
    `include "LTSSM1_seq_item.sv"
    `include "LTSSM2_seq_item.sv"
    `include "PIPE_seq_item.sv"
    `include "TX_Master_seq_item.sv"// CHANGE 

    `include "Reset_LTSSM1_seq.sv"
    `include "Reset_LTSSM2_seq.sv"
    `include "LinkUp1_seq.sv"
    `include "LinkUp2_seq.sv"
    `include "TLP_Seq_TX_MASTER_D.sv"
    `include "TLP_Seq_TX_MASTER_U.sv"
    `include "DLLP_Seq_TX_MASTER_D.sv"
    `include "DLLP_Seq_TX_MASTER_U.sv"
    `include "DLLP_TLP_Seq_TX_MASTER_D.sv"
    `include "DLLP_TLP_Seq_TX_MASTER_U.sv"


    `include "RX_Slave_Config.sv"
    `include "TX_Slave_Config.sv"
    `include "LTSSM1_Config.sv"
    `include "LTSSM2_Config.sv"
    `include "TX_Master_Config.sv"
    `include "RX_Passive_Config.sv"

    `include "RX_Slave_D_Monitor.sv"
    `include "RX_Slave_D_Driver.sv"
    `include "RX_Slave_D_Agent.sv"
    `include "RX_Slave_U_Monitor.sv"
    `include "RX_Slave_U_Driver.sv"
    `include "RX_Slave_U_Agent.sv"
    

    `include "TX_Slave_D_Monitor.sv"
    `include "TX_Slave_D_Agent.sv"
    `include "TX_Slave_U_Monitor.sv"
    `include "TX_Slave_U_Agent.sv"
    
    `include "TX_Master_D_Sequencer.sv"
    `include "TX_Master_D_Driver.sv"
    `include "TX_Master_D_Agent.sv"

    `include "TX_Master_U_Sequencer.sv"
    `include "TX_Master_U_Driver.sv"
    `include "TX_Master_U_Agent.sv"

    
    `include "RX_Passive_D_Monitor.sv"
    `include "RX_Passive_D_Agent.sv"

    `include "RX_Passive_U_Monitor.sv"
    `include "RX_Passive_U_Agent.sv"

    

    

    `include "LTSSM1_D_Driver.sv"
   // `include "LTSSM1_D_Monitor.sv"
    `include "LTSSM1_D_Sequencer.sv"
    `include "LTSSM1_D_Agent.sv"
    
    
    `include "LTSSM1_U_Driver.sv"
    //`include "LTSSM1_U_Monitor.sv"
    `include "LTSSM1_U_Sequencer.sv"
    `include "LTSSM1_U_Agent.sv"



    `include "LTSSM2_D_Driver.sv"
    `include "LTSSM2_D_Monitor.sv"
    `include "LTSSM2_D_Sequencer.sv"
    `include "LTSSM2_D_Agent.sv"
    
    
    `include "LTSSM2_U_Driver.sv"
    `include "LTSSM2_U_Monitor.sv"
    `include "LTSSM2_U_Sequencer.sv"
    `include "LTSSM2_U_Agent.sv"

    `include "LinkUp1_vseq.sv"
    `include "LinkUp2_vseq.sv"

    `include "TLP_vSeq_TX_MASTER.sv"
    `include "DLLP_vSeq_TX_MASTER.sv"
    `include "DLLP_TLP_vSeq_TX_MASTER.sv"

    `include "Adapter.sv"

    `include "PCIe_Env.sv"

    `include "PCIe_Test.sv"
    
    
endpackage
