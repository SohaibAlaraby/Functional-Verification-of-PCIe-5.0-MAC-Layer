class RX_Slave_U_Monitor  extends uvm_monitor;
  
`uvm_component_utils(RX_Slave_U_Monitor)


virtual PIPE_if PIPE_vif_h; 

uvm_analysis_port #(PIPE_seq_item) send_ap;


extern function new(string name="RX_Slave_U_Monitor",uvm_component parent);
extern function void build_phase(uvm_phase phase);
extern function void connect_phase(uvm_phase phase);
extern task run_phase(uvm_phase phase);

    

endclass







function RX_Slave_U_Monitor::new(string name="RX_Slave_U_Monitor",uvm_component parent);
  
        super.new(name,parent);

        
endfunction 




function void RX_Slave_U_Monitor::build_phase(uvm_phase phase);
  
        super.build_phase(phase);
        `uvm_info(get_type_name() ," in monitor build_phase ",UVM_HIGH)
       
        send_ap = new("send_ap",this);
                
endfunction




function void RX_Slave_U_Monitor::connect_phase(uvm_phase phase);
  
        super.connect_phase(phase);
        `uvm_info(get_type_name() ," in monitor connect_phase ",UVM_HIGH)
        
endfunction
   
   
   
   
    
task RX_Slave_U_Monitor::run_phase(uvm_phase phase);
        super.run_phase(phase);
        `uvm_info(get_type_name() ," in monitor run_phase ",UVM_HIGH)
        //forever begin
         
       // end
endtask
    