`ifndef MAXPIPEWIDTH
`define MAXPIPEWIDTH 32;
`endif

`ifndef MAXPIPEWIDTH
`define LANESNUMBER 16;
`endif