

`ifndef MAXPIPEWIDTH
   `define MAXPIPEWIDTH 32
`endif

`ifndef LANESNUMBER
   `define LANESNUMBER 16
`endif

`define MAX_GEN_PCIE_D 1 
`define MAX_GEN_PCIE_U 1 