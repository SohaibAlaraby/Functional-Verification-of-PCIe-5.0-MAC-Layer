package PCIe_pkg;
    import uvm_pkg::*;
    
    `include "uvm_macros.svh"
    `include "Defines.sv"
    `include "PCIe_Seq_Item.sv"
    `include "PCIe_Sequence_AUM.sv"
    `include "PCIe_Sequence_ADM.sv"
    `include "PCIe_Sequencer_AUM.sv"
    `include "PCIe_Sequencer_ADM.sv"

    `include "PCIe_Driver_AUM.sv"
    `include "PCIe_Driver_ADM.sv"
    `include "PCIe_Driver_AUS2.sv"
    `include "PCIe_Driver_ADS2.sv"
    
    `include "PCIe_Monitor_ADL1.sv"
    `include "PCIe_Monitor_ADL2.sv"
    `include "PCIe_Monitor_ADM.sv"
    `include "PCIe_Monitor_ADS1.sv"
    `include "PCIe_Monitor_ADS2.sv"
    `include "PCIe_Monitor_ADS3.sv"
    `include "PCIe_Monitor_AUL1.sv"
    `include "PCIe_Monitor_AUL2.sv"
    `include "PCIe_Monitor_AUM.sv"
    `include "PCIe_Monitor_AUS1.sv"
    `include "PCIe_Monitor_AUS2.sv"
    `include "PCIe_Monitor_AUS3.sv"

    `include "PCIe_CoverageCollector_D.sv"
    `include "PCIe_CoverageCollector_U.sv"

    `include "PCIe_ScoreboardD.sv"
    `include "PCIe_ScoreboardU.sv"

    `include "PCIe_AgentD_LTSSM1.sv"
    `include "PCIe_AgentD_LTSSM2.sv"
    `include "PCIe_AgentD_Master.sv"
    `include "PCIe_AgentD_Slave1.sv"
    `include "PCIe_AgentD_Slave2.sv"
    `include "PCIe_AgentD_Slave3.sv"
    `include "PCIe_AgentU_LTSSM1.sv"
    `include "PCIe_AgentU_LTSSM2.sv"
    `include "PCIe_AgentU_Master.sv"
    `include "PCIe_AgentU_Slave1.sv"
    `include "PCIe_AgentU_Slave2.sv"
    `include "PCIe_AgentU_Slave3.sv"

    `include "PCIe_Env.sv"

    `include "PCIe_Test0.sv"
endpackage