class TX_Slave_U_Monitor extends uvm_monitor;
  


`uvm_component_utils(TX_Slave_U_Monitor)
    

virtual PIPE_if      PIPE_vif_h;
 
uvm_analysis_port #(PIPE_TX_seq_item_h) send_ap1;
uvm_analysis_port #(PIPE_TX_seq_item_h) send_ap2;

    
extern function new(string name = "TX_Slave_U_Monitor",uvm_component parent);
extern function void build_phase (uvm_phase phase);
extern function void connect_phase (uvm_phase phase);
extern task run_phase(uvm_phase phase);
extern task Pass_PIPE_TX_Signals ();



endclass






function TX_Slave_U_Monitor::new(string name = "TX_Slave_U_Monitor",uvm_component parent);
        super.new(name , parent);
        `uvm_info(get_type_name() ," in constructor of driver ",UVM_HIGH)
endfunction 



function void TX_Slave_U_Monitor::build_phase (uvm_phase phase);
  
        super.build_phase(phase);
        
        `uvm_info(get_type_name() ," in build_phase of driver ",UVM_LOW)
        
        send_ap1 = new("send_ap1",this);
        send_ap2 = new("send_ap2",this);   
             
endfunction: build_phase



function void TX_Slave_U_Monitor::connect_phase (uvm_phase phase);
        super.connect_phase(phase);
        `uvm_info(get_type_name() ," in connect_phase of driver ",UVM_LOW)
endfunction: connect_phase





task TX_Slave_U_Monitor::run_phase(uvm_phase phase);
  
        super.run_phase(phase);
        `uvm_info(get_type_name() ," in run_phase of driver ",UVM_LOW)
      
        fork
        
              Pass_PIPE_TX_Signals();
        
        join
        
endtask: run_phase





task TX_Slave_U_Monitor::Pass_PIPE_TX_Signals();
  
  forever begin
    
     PIPE_TX_seq_item  PIPE_TX_seq_item_h;         
     PIPE_TX_seq_item_h = PIPE_TX_seq_item::type_id::create("PIPE_TX_seq_item_h"); 
     
     @(posedge PIPE_vif_h.CLK)   
  
     PIPE_TX_seq_item_h.TxData                  = PIPE_vif_h.TxData;
     PIPE_TX_seq_item_h.TxDataValid             = PIPE_vif_h.TxDataValid;
     PIPE_TX_seq_item_h.TxElecIdle              = PIPE_vif_h.TxElecIdle;
     PIPE_TX_seq_item_h.TxStartBlock            = PIPE_vif_h.TxStartBlock;
     PIPE_TX_seq_item_h.TxDataK                 = PIPE_vif_h.TxDataK;
     PIPE_TX_seq_item_h.TxSyncHeader            = PIPE_vif_h.TxSyncHeader;
     PIPE_TX_seq_item_h.TxDetectRx_Loopback     = PIPE_vif_h.TxDetectRx_Loopback;
     
     send_ap1.write(PIPE_TX_seq_item_h);
    
   end
  

endtask