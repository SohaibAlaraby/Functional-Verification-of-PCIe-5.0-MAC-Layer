

`ifndef MAXPIPEWIDTH
   `define MAXPIPEWIDTH 32
`endif

`ifndef LANESNUMBER
   `define LANESNUMBER 16
`endif